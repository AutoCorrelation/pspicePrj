** Profile: "SCHEMATIC1-p176"  [ c:\users\user\desktop\codespace\pspiceprj\exp6_1-PSpiceFiles\SCHEMATIC1\p176.sim ] 

** Creating circuit file "p176.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.OP
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
